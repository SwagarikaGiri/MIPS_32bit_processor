 module register_file (clk,rst,r_wr_en,r_reg1,r_reg2,w_reg,w_data,r1_data,r2_data) ;
 
      input clk;
	  input rst;
      input r_wr_en;
	  input [4:0] r_reg1;
	  input [4:0]  r_reg2;
	  input [4:0] w_reg;
	  output [31:0] r1_data;
	  output [31:0] r2_data;
	  input [31:0] w_data;
      reg [31:0] memdata [31:0];
      
   
      
     initial
        begin
        

         memdata[0] = 32'b00000000001000100001100000100000;
         memdata[1] = 32'b00000000001000100001100000100010;
		 memdata[2] = 32'b00000000001000100001100000100011;
		 memdata[3] = 32'b00000000001000100001100000100101;
		 memdata[4] = 32'b10000000001000100001100000100000;
		 memdata[5] = 32'b00000000001000100001100000100000;
         memdata[6] = 32'b00000000001000100001100000100010;
		 memdata[7] = 32'b00000000001000100001100000100100;
		 memdata[8] = 32'b00000000001000100001100000100101;
		 memdata[9] = 32'b10000000001000100001100000100000;
		memdata[10] = 32'b00000000001000100001100000100000;
        memdata[11] = 32'b00000000001000100001100000100010;
		memdata[12] = 32'b00000000001000100001100000100100;
		memdata[13] = 32'b00000000001000100001100000100101;
		memdata[14] = 32'b10000000001000100001100000100000;
		memdata[15] = 32'b00000000001000100001100000100000;
        memdata[16] = 32'b00000000001000100001100000100010;
		memdata[17] = 32'b00000000001000100001100000100100;
		memdata[18] = 32'b00000000001000100001100000100101;
		memdata[19] = 32'b10000000001000100001100000100000;
		memdata[20] = 32'b00000000001000100001100000100000;
        memdata[21] = 32'b00000000001000100001100000100010;
		memdata[22] = 32'b00000000001000100001100000100100;
		memdata[23] = 32'b00000000001000100001100000100101;
		memdata[24] = 32'b10000000001000100001100000100000;
		memdata[25] = 32'b00000000001000100001100000100000;
        memdata[26] = 32'b00000000001000100001100000100010;
		memdata[27] = 32'b00000000001000100001100000100100;
		memdata[28] = 32'b00000000001000100001100000100101;
		memdata[29] = 32'b10000000001000100001100000100000;
		memdata[30] = 32'b00000000001000100001100000100000;
        memdata[31] = 32'b00000000001000100001100000100010;
  end
      assign  r1_data=memdata[r_reg1]; 
	  assign  r2_data=memdata[r_reg2];
	     /* always
	    begin
		  if(r_wr_en ==1'b1)
		   begin 
		    memdata[w_reg] == w_data;
		  end
		end  */
		
	  
  endmodule
  